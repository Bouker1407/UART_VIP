interface uart_if();

  logic TX;
  logic RX;
  
endinterface
